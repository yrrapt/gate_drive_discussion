********************************************************************************
* UnitedSiC G3 1200V-140mohm SiC JFET Spice Circuit Model v3.1
* Copyright 2018 United Silicon Carbide, Inc.
* This is a PRELIMINARY Spice Model of UF3N120140Z
*
*
* The model does not include all possible conditions and effects,
* in particular it doesn't include:
*	Self heating
*	leakage current in blocking state
*	Drain to source breakdown is notional only
*
********************************************************************************


*** UF3N120140Z ***
.subckt UF3N120140Z nd ng ns
*#ASSOC Category="N-Channel JFET" Symbol=njfet
xj1	nd	ng	ns	jfet_G3_1200V_Ron params: Ron=140m Rgoff=1.6 Rgon=1.6
.ends

*** 1200V JFETs ***
.subckt jfet_G3_1200V_Ron d g s params: Ron=0 Rgon=0 Rgoff=0
.param Ron1={Ron}
.param Rgon1={Rgon}
.param Rgoff1={Rgoff}
.param a= {75m / {Ron1}}
X1 di gi s jfet_G3_1200V params: ascale={a}
XCgs gi s Cgs_1200V params: acgs={a}
XCgd gi di Cgd_1200V params: acgd={a}
Cgdex gi di {25p * {a} }
Cgsex gi s {0.2n * {a} }
Rd d di Rtemp {58.2m/{a}}
.MODEL Rtemp RES (TC1=3.93e-3, TC2=4.79e-5)
GRg g gi value={if(v(g,gi)>0,v(g,gi)/{Rgon1},v(g,gi)/{Rgoff1})}
.ends jfet_G3_1200V_Ron

*** Shared Subcircuit for 1200V JFETs ***
.subckt jfet_G3_1200V d g s Params: ascale=0
.param Fc1=0.5
.param Pb1=3.25
.param M1=0.5
.param Vd0=800

.param gos={0.0178*{ascale}}
.param gfs={43*{ascale}}
.param f=1.453
.param vth=-11.5

.param cgs1=0.594n
.param cgd1=0.0318n

.param bt={({f}*{gfs}+2*{gos}*{Vd0}/{vth})/2/(-{vth})}
.param lamd={1*{gos}/{bt}/{vth}/{vth}}
.param cgs0={pwr((1+30/{Pb1}),{M1})*{cgs1}}
.param cgd0={pwr((1+{Vd0}/{Pb1}),{M1})*{cgd1}}

J1 d g s jfet_1200
Dgs g s Dgs_iv
Dgd g d Dgd_iv
Rgs  g s 1Meg
Rgd  g d 10Meg

.MODEL jfet_1200 NJF(
+ Beta={bt} BetaTce=0 Vto={vth} VtoTc=0  lambda={lamd}
+ Is=1e-60
+ Cgs={{cgs0}*{ascale}} Cgd={{cgd0}*{ascale}} Fc={Fc1} Pb={Pb1}
+ M={M1})

.MODEL Dgs_iv D (CJO=0 BV=40 IS=1e-50 ISR=1e-50 Eg=3.5 Rs=0)
.MODEL Dgd_iv D (CJO=0 BV=1500 IS=1e-50 ISR=1e-50 Eg=3.5 Rs={9.62m/{ascale}})
.ends jfet_G3_1200V

* Cgs network
.subckt Cgs_1200V g s params: acgs=0
.param c0=1n
.param vsgmin=-2
.param vsgmax=15
.param a1={0.8n*{acgs}}
.param b1=1
.func Qgs1(u) {- {a1} / {b1} *(exp(- {b1} *u)-1)}


.param a2={0.7n*{acgs}}
.param b2=0.75
.param c2=9.5


.func Qgs2(u)
+	{if(abs(u)<{vsgmax},
+	{a2}*u + {a2}*(-{b2})*log(cosh((u-{c2})/-{b2}))
+	-{a2}*(-{b2})*log(cosh(-{c2}/-{b2})),
+	{a2}*{vsgmax} + {a2}*(-{b2})*log(cosh(({vsgmax}-{c2})/-{b2}))
+	-{a2}*(-{b2})*log(cosh(-{c2}/-{b2})))}


E1 s m1 value={v(s,g)-Qgs1(v(s,g))/{c0}}
C01 m1 g {c0}
E2 s m2 value={v(s,g)-Qgs2(limit(v(s,g),-{vsgmax},{vsgmax}))/{c0}}
C02 m2 g {c0}

.ends Cgs_1200V

* Cgd network
.subckt Cgd_1200V g d params:acgd=0

.param c0=1n

.param a1={0.3n*{acgd}}
.param b1=0.9
.param c1=20
.param vdgmax1=30

.func Qgd1(u)
+	{if(abs(u)<{vdgmax1},
+	{a1}*u + {a1}*(-{b1})*log(cosh((u-{c1})/-{b1}))
+	-{a1}*(-{b1})*log(cosh(-{c1}/-{b1})),
+	{a1}*{vdgmax1} + {a1}*(-{b1})*log(cosh(({vdgmax1}-{c1})/-{b1}))
+	-{a1}*(-{b1})*log(cosh(-{c1}/-{b1})))}

.param a2={0*{acgd}}
.param b2=0.5
.param c2=9.5
.param vdgmax2=15

.func Qgd2(u)
+	{if(abs(u)<{vdgmax2},
+	(-1)*({a2}*u + {a2}*(-{b2})*log(cosh((u-{c2})/-{b2}))
+	-{a2}*(-{b2})*log(cosh(-{c2}/-{b2}))),
+	(-1)*({a2}*{vdgmax2} + {a2}*(-{b2})*log(cosh(({vdgmax2}-{c2})/-{b2}))
+	-{a2}*(-{b2})*log(cosh(-{c2}/-{b2}))))}

E1 d m1 value={v(d,g)-Qgd1(limit(v(d,g),-{vdgmax1},+{vdgmax1}))/{c0}}
C01 m1 g {c0}
E2 d m2 value={v(d,g)-Qgd2(limit(v(d,g),-{vdgmax2},+{vdgmax2}))/{c0}}
C02 m2 g {c0}

.ends Cgd_1200V

*** End of File ***
